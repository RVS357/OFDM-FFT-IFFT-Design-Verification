interface ofdm_intf(input Clk, input Reset);

 logic Pushin;
 logic FirstData;
 logic signed [16:0] DinR;
 logic signed [16:0] DinI;
 logic PushOut;
 logic [47:0] DataOut;
  
  //modport

endinterface
